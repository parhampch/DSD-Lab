module Booth(
    input [4:0] a,
    input [4:0] b,
    input clk,
    input rst,
    output [9:0] c,
    output done);


    
endmodule